`timescale 1 ns / 1 ps

module XNORARRAY_b0 (
        lut_out_63_V_write,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63);

parameter    ap_const_lv288_0_0 = 288'h3F51F7D81DD70FB9DED197B8439087C4765E9A1B77D73A96E915C7D3751FBCAE799198B8;
parameter    ap_const_lv288_0_1 = 288'hDD99E4D6CF19E4DA322FE802B10F8D1027DEAE5232FFE8B9348E8938260A9EAD2E1EB9B0;
parameter    ap_const_lv288_0_2 = 288'hC955BD98C95536C8F9136C4A67AD9817F73DB74B5931E01B90A61D4401C5CC2C046D4880;
parameter    ap_const_lv288_0_3 = 288'h8F1C88D123FE2A0FB27E29200158844097B9DEFBAFFFBA7B1190B0C10119B19B272FBE97;
parameter    ap_const_lv288_0_4 = 288'h778289756E179920237FEA2820418912058BC83038FF892B0A52C8A9026649993C3F8C36;
parameter    ap_const_lv288_0_5 = 288'hFDBFBE5FFBBF3757B3BF3F7FB4EF5E5EAFEA7E469BFF3F5A7F819E7AFF91F67CFFB7B64A;
parameter    ap_const_lv288_0_6 = 288'h75E66820DDC9BD746D18E7DF75E7E932B5EE23746F98A68EF093B830ED25FB7FCD90B7CF;
parameter    ap_const_lv288_0_7 = 288'h7D5F4EFF742E5E272DAB5E2E599B8AD8CE9A0EFA99C116DE745D46AA6C7A7EA4683A25C2;
parameter    ap_const_lv288_0_8 = 288'hD9C9C7D659B9E4D12B7A242B7022C942C100A91D07F8B69BD4E61970C4ACCB4C4589B65F;
parameter    ap_const_lv288_0_9 = 288'hF2D176CED1D8751AD9B975D77F73F07FD9E15B7AF9A97757F7A9E0C7D80543079B29665F;
parameter    ap_const_lv288_0_10 = 288'hFC83B916D38BA88622AF680372ABA052D1DDE1E3063D6C8F80EFB92A00E6A961027E6F26;
parameter    ap_const_lv288_0_11 = 288'hD91F4900A44C68A7AFE66232B1480940216DE4A38EF7F6B7390A49523D4E60D9ED76E23;
parameter    ap_const_lv288_0_12 = 288'h2684086B34DE9D792A9C5D5ACAA7B2F71EA2839A67E216195E63B6A98E68F98887E2F2B;
parameter    ap_const_lv288_0_13 = 288'h660E1005010E0805651C7B2A058F002DA45E7E91AE762B8C5A8F004773E715036EE3A39;
parameter    ap_const_lv288_0_14 = 288'h6A68C2AF3468C3B632ACC175BEFE66AA7A6074BC82EE2551573C936B9E6B674E8E7E677B;
parameter    ap_const_lv288_0_15 = 288'hB58E68100501981459191BC0A70D588B1D085A0DD45819181D545D998CD45435C4D8126;
parameter    ap_const_lv288_0_16 = 288'h7547883027CB32BE6218722E750990BC16F170BC88F2742C6A5B5ABA5870728882B4734B;
parameter    ap_const_lv288_0_17 = 288'h7987DF343F81CCB27853CC9A76036C6D924DF79F7987C881326B0F3B1E372905B8260D07;
parameter    ap_const_lv288_0_18 = 288'h8220704E842851870028400787EC736FC729126D6F6EC57DDDE5334B5CEF3B38CEFF4331;
parameter    ap_const_lv288_0_19 = 288'h80003C544C17B888F997BA882778F6573604E8A63B97B893A88ABE79A5EEE93A3F97FC98;
parameter    ap_const_lv288_0_20 = 288'h76229885D789919D99C5DCDAE6CBD8ADC76BB5EB3AF6C468244ABA212E78A6AA2A560CA0;
parameter    ap_const_lv288_0_21 = 288'hCBD596D9A36E5A2C3DF71BE8CF720E0A7FE25E7CBFFF1B50673952AA7F3BDAFD7FB7BBDC;
parameter    ap_const_lv288_0_22 = 288'h608608058A1D3892F7955BED8003894ADD5CD2927FDE93EB84E7A84791F6EF4BD5E9767D;
parameter    ap_const_lv288_0_23 = 288'h3FFD777E74BC27395FC1D7FDBFB2D67A10B40FE5212495ADF5E0376ABFE966D7F360577B;
parameter    ap_const_lv288_0_24 = 288'h895DC7CB8A6D420BA26E690382CC86D8FFEB5A7FA6EE2F71026C318DCA2F4B0D8E7E6FC7;
parameter    ap_const_lv288_0_25 = 288'h122E7A0F32AE097786440954862FBB6BB9B07E5F0E7F2F75D7ECBB78ADAEAFEB8E5E3F43;
parameter    ap_const_lv288_0_26 = 288'h79D5BD910B15BCC8F991B28B4B194096465850E67F01D0962A7846AB7C50523335AA4034;
parameter    ap_const_lv288_0_27 = 288'h59D8959040500985440040A44A1D3BB06812AAA96E50A9AF4B5C86E3775686887050CC28;
parameter    ap_const_lv288_0_28 = 288'hC60608806002D8803807DA8206DA7B65F0C259247982C8823A6A6B2C20226BB120C69DDD;
parameter    ap_const_lv288_0_29 = 288'h8217198C0013184D08115A892E1D06E624552792AD1110B0F5B66FC3F2D22EF3F598F775;
parameter    ap_const_lv288_0_30 = 288'hB463B86475BBE85BBFEF3A7298E46141906A71479ABA47528664C98483E3521DCA3B574A;
parameter    ap_const_lv288_0_31 = 288'h1FF9F6FFDE39F7D9CF1087DD5DEDE29E9EE1D41BDD91B157C0FC21C09CED5C0CD80150D4;
parameter    ap_const_lv288_0_32 = 288'h9A87AC5089C53752FFD176D86303E846DFAE7A7873B850F9CA4F0A33862EBBA5B1E55468;
parameter    ap_const_lv288_0_33 = 288'h908F8993D7D7AA9E82F48918640A8AA286DBA6AA48F7CD20615C98A2675CA0A26856A1A0;
parameter    ap_const_lv288_0_34 = 288'h59FDC3B925B8C6331E6075FD744B9FBECA5B2F9E47FC6276751B1EAE6B52560EDF5D67DC;
parameter    ap_const_lv288_0_35 = 288'hE4F6A949E7BEABED863E2A21661398284399B6CA6C54FE277813AC270191945651D4D246;
parameter    ap_const_lv288_0_36 = 288'h5959C7D9006D40B7262A783710654050413D5854D7A832FD70E78BBD50465EE58DE8720F;
parameter    ap_const_lv288_0_37 = 288'hA6A628478E33B94DD1BFC84185A7397B6FC485E080669FD300EE690820E68D733CBA6895;
parameter    ap_const_lv288_0_38 = 288'h27B7187DAF96BF7DDF971AF8AF9BAE5DAE9FA4DD1D5318F0ED929FF2ABF1E461B5C61930;
parameter    ap_const_lv288_0_39 = 288'hC27073EB90C8555785287567CF3753DFD9E3533CC5E8714717ED57731AE74FFED1ED7255;
parameter    ap_const_lv288_0_40 = 288'hE7CC6EF3E6C47E7066C612618DEA6481E4A2F978A5F6B2451BD84DF5F7FA2CAC21EA287;
parameter    ap_const_lv288_0_41 = 288'h78578F392D8F0AB82C17380A7F1F4CFBA43C12668518F00FFA1B0ECB98740F16987117CE;
parameter    ap_const_lv288_0_42 = 288'h7549C492791DC4B04C01C493329A58BFFA02A81490404D343CF25ECC087E6B39464E0BA5;
parameter    ap_const_lv288_0_43 = 288'h5941E59055D584BD7F98E67B12406120140488D1FD11F29F1265413080C81960C489D5CE;
parameter    ap_const_lv288_0_44 = 288'h7581E6B02964E4DCD819668B7331F094407668588A1C67437F39A0EE6C7624FD8E4C73A9;
parameter    ap_const_lv288_0_45 = 288'h8678766FF6E2566AB0E640550FE8766AFF1BBBDDBFB70BD8A4EC276BAECBBE382EEF1A38;
parameter    ap_const_lv288_0_46 = 288'h7C8F9F307B8FAEDEAE7F2A23655E8CE0C171F70737B9503898DD2DD9514110F884A1D1FA;
parameter    ap_const_lv288_0_47 = 288'hB26279227BA96851D359F3F7BEEA2963794BBDD7F011F49F84A27B47356CE814F930C4CB;
parameter    ap_const_lv288_0_48 = 288'h35D32FB06CB03C3C799195DC7911305858141148FEB3C4D37E1B46D9083E45D99F2D6635;
parameter    ap_const_lv288_0_49 = 288'h8666992886EA99A405E489F582C23BA871C0572159D8352ED354B5875BF1327EF99194FE;
parameter    ap_const_lv288_0_50 = 288'hF9F48DD81AD78DD3261F09A199D62D16262E6F7377187AB79C4F1BB0B5A9F8FCF599F4DF;
parameter    ap_const_lv288_0_51 = 288'h82F071E991F841E7A52C64278DC6A7DB99459F508588A736046F4B356EC68AA8D0FD1BCC;
parameter    ap_const_lv288_0_52 = 288'h362A88A017F9A1BF826C6D23201AA8A700EA27AA6A74EF630222C9AA41368ECAC87C0703;
parameter    ap_const_lv288_0_53 = 288'h24E8F0069679F3BA75D9D7DFA4AC5900C609F937BD9197DA80A4116537AD995135D9B7DE;
parameter    ap_const_lv288_0_54 = 288'h424031244754A9882012A8005041A091541EA590A5D0AC1317E5A0DC07A8A0EE1CE1D462;
parameter    ap_const_lv288_0_55 = 288'h3FB2762EB1B8E9F33FE8E57528A1B60A9EA057DD3BF8AF94E72D936EEFF9F6FF07D82658;
parameter    ap_const_lv288_0_56 = 288'hA4071D84C90598C0AB17AE8A870F891DCE0DB1A2652FC88A02C749144044492048A64826;
parameter    ap_const_lv288_0_57 = 288'h753669F162B66547066E6B2788570D90C809D38B827AC6015D8FF2B11D2EE7971E176034;
parameter    ap_const_lv288_0_58 = 288'h7FEFEE7E79BE7E187BD73EDC7F2BEE7F7B9BFE3D7F367C9A3E382ED43F3AB8C47B373AB9;
parameter    ap_const_lv288_0_59 = 288'h9DFF47BB2E4F4A82765789909C7E4F22FCB1586535C79930075C5BAA75D08F9737C3A933;
parameter    ap_const_lv288_0_60 = 288'hA0B23C6DBE7B3677B1AE3D7D8C3A2E4FAD6977DFFBBE3B7DADEE7F7EECEA5E49ABFE3E7C;
parameter    ap_const_lv288_0_61 = 288'h7D81F7B07B81E6885A5D66F279D4A49498162C0050686603795D84D98A765CA890665A29;
parameter    ap_const_lv288_0_62 = 288'h82A719598B3F1B4DB9B61A5DCE673A4FEFEC3A64D7A33CD8674F8AA36701F2A871F35AE8;
parameter    ap_const_lv288_0_63 = 288'h19BCA65A89DDC74B7E196E3399B0755ABA082F477E1BBE07BD31F7DDF3BD1657F91FA44D;


input  [287:0] lut_out_63_V_write;
output  [287:0] ap_return_0;
output  [287:0] ap_return_1;
output  [287:0] ap_return_2;
output  [287:0] ap_return_3;
output  [287:0] ap_return_4;
output  [287:0] ap_return_5;
output  [287:0] ap_return_6;
output  [287:0] ap_return_7;
output  [287:0] ap_return_8;
output  [287:0] ap_return_9;
output  [287:0] ap_return_10;
output  [287:0] ap_return_11;
output  [287:0] ap_return_12;
output  [287:0] ap_return_13;
output  [287:0] ap_return_14;
output  [287:0] ap_return_15;
output  [287:0] ap_return_16;
output  [287:0] ap_return_17;
output  [287:0] ap_return_18;
output  [287:0] ap_return_19;
output  [287:0] ap_return_20;
output  [287:0] ap_return_21;
output  [287:0] ap_return_22;
output  [287:0] ap_return_23;
output  [287:0] ap_return_24;
output  [287:0] ap_return_25;
output  [287:0] ap_return_26;
output  [287:0] ap_return_27;
output  [287:0] ap_return_28;
output  [287:0] ap_return_29;
output  [287:0] ap_return_30;
output  [287:0] ap_return_31;
output  [287:0] ap_return_32;
output  [287:0] ap_return_33;
output  [287:0] ap_return_34;
output  [287:0] ap_return_35;
output  [287:0] ap_return_36;
output  [287:0] ap_return_37;
output  [287:0] ap_return_38;
output  [287:0] ap_return_39;
output  [287:0] ap_return_40;
output  [287:0] ap_return_41;
output  [287:0] ap_return_42;
output  [287:0] ap_return_43;
output  [287:0] ap_return_44;
output  [287:0] ap_return_45;
output  [287:0] ap_return_46;
output  [287:0] ap_return_47;
output  [287:0] ap_return_48;
output  [287:0] ap_return_49;
output  [287:0] ap_return_50;
output  [287:0] ap_return_51;
output  [287:0] ap_return_52;
output  [287:0] ap_return_53;
output  [287:0] ap_return_54;
output  [287:0] ap_return_55;
output  [287:0] ap_return_56;
output  [287:0] ap_return_57;
output  [287:0] ap_return_58;
output  [287:0] ap_return_59;
output  [287:0] ap_return_60;
output  [287:0] ap_return_61;
output  [287:0] ap_return_62;
output  [287:0] ap_return_63;
assign ap_return_0 = ~(ap_const_lv288_0_0 ^ lut_out_63_V_write);
assign ap_return_1 = ~(ap_const_lv288_0_1 ^ lut_out_63_V_write);
assign ap_return_2 = ~(ap_const_lv288_0_2 ^ lut_out_63_V_write);
assign ap_return_3 = ~(ap_const_lv288_0_3 ^ lut_out_63_V_write);
assign ap_return_4 = ~(ap_const_lv288_0_4 ^ lut_out_63_V_write);
assign ap_return_5 = ~(ap_const_lv288_0_5 ^ lut_out_63_V_write);
assign ap_return_6 = ~(ap_const_lv288_0_6 ^ lut_out_63_V_write);
assign ap_return_7 = ~(ap_const_lv288_0_7 ^ lut_out_63_V_write);
assign ap_return_8 = ~(ap_const_lv288_0_8 ^ lut_out_63_V_write);
assign ap_return_9 = ~(ap_const_lv288_0_9 ^ lut_out_63_V_write);
assign ap_return_10 = ~(ap_const_lv288_0_10 ^ lut_out_63_V_write);
assign ap_return_11 = ~(ap_const_lv288_0_11 ^ lut_out_63_V_write);
assign ap_return_12 = ~(ap_const_lv288_0_12 ^ lut_out_63_V_write);
assign ap_return_13 = ~(ap_const_lv288_0_13 ^ lut_out_63_V_write);
assign ap_return_14 = ~(ap_const_lv288_0_14 ^ lut_out_63_V_write);
assign ap_return_15 = ~(ap_const_lv288_0_15 ^ lut_out_63_V_write);
assign ap_return_16 = ~(ap_const_lv288_0_16 ^ lut_out_63_V_write);
assign ap_return_17 = ~(ap_const_lv288_0_17 ^ lut_out_63_V_write);
assign ap_return_18 = ~(ap_const_lv288_0_18 ^ lut_out_63_V_write);
assign ap_return_19 = ~(ap_const_lv288_0_19 ^ lut_out_63_V_write);
assign ap_return_20 = ~(ap_const_lv288_0_20 ^ lut_out_63_V_write);
assign ap_return_21 = ~(ap_const_lv288_0_21 ^ lut_out_63_V_write);
assign ap_return_22 = ~(ap_const_lv288_0_22 ^ lut_out_63_V_write);
assign ap_return_23 = ~(ap_const_lv288_0_23 ^ lut_out_63_V_write);
assign ap_return_24 = ~(ap_const_lv288_0_24 ^ lut_out_63_V_write);
assign ap_return_25 = ~(ap_const_lv288_0_25 ^ lut_out_63_V_write);
assign ap_return_26 = ~(ap_const_lv288_0_26 ^ lut_out_63_V_write);
assign ap_return_27 = ~(ap_const_lv288_0_27 ^ lut_out_63_V_write);
assign ap_return_28 = ~(ap_const_lv288_0_28 ^ lut_out_63_V_write);
assign ap_return_29 = ~(ap_const_lv288_0_29 ^ lut_out_63_V_write);
assign ap_return_30 = ~(ap_const_lv288_0_30 ^ lut_out_63_V_write);
assign ap_return_31 = ~(ap_const_lv288_0_31 ^ lut_out_63_V_write);
assign ap_return_32 = ~(ap_const_lv288_0_32 ^ lut_out_63_V_write);
assign ap_return_33 = ~(ap_const_lv288_0_33 ^ lut_out_63_V_write);
assign ap_return_34 = ~(ap_const_lv288_0_34 ^ lut_out_63_V_write);
assign ap_return_35 = ~(ap_const_lv288_0_35 ^ lut_out_63_V_write);
assign ap_return_36 = ~(ap_const_lv288_0_36 ^ lut_out_63_V_write);
assign ap_return_37 = ~(ap_const_lv288_0_37 ^ lut_out_63_V_write);
assign ap_return_38 = ~(ap_const_lv288_0_38 ^ lut_out_63_V_write);
assign ap_return_39 = ~(ap_const_lv288_0_39 ^ lut_out_63_V_write);
assign ap_return_40 = ~(ap_const_lv288_0_40 ^ lut_out_63_V_write);
assign ap_return_41 = ~(ap_const_lv288_0_41 ^ lut_out_63_V_write);
assign ap_return_42 = ~(ap_const_lv288_0_42 ^ lut_out_63_V_write);
assign ap_return_43 = ~(ap_const_lv288_0_43 ^ lut_out_63_V_write);
assign ap_return_44 = ~(ap_const_lv288_0_44 ^ lut_out_63_V_write);
assign ap_return_45 = ~(ap_const_lv288_0_45 ^ lut_out_63_V_write);
assign ap_return_46 = ~(ap_const_lv288_0_46 ^ lut_out_63_V_write);
assign ap_return_47 = ~(ap_const_lv288_0_47 ^ lut_out_63_V_write);
assign ap_return_48 = ~(ap_const_lv288_0_48 ^ lut_out_63_V_write);
assign ap_return_49 = ~(ap_const_lv288_0_49 ^ lut_out_63_V_write);
assign ap_return_50 = ~(ap_const_lv288_0_50 ^ lut_out_63_V_write);
assign ap_return_51 = ~(ap_const_lv288_0_51 ^ lut_out_63_V_write);
assign ap_return_52 = ~(ap_const_lv288_0_52 ^ lut_out_63_V_write);
assign ap_return_53 = ~(ap_const_lv288_0_53 ^ lut_out_63_V_write);
assign ap_return_54 = ~(ap_const_lv288_0_54 ^ lut_out_63_V_write);
assign ap_return_55 = ~(ap_const_lv288_0_55 ^ lut_out_63_V_write);
assign ap_return_56 = ~(ap_const_lv288_0_56 ^ lut_out_63_V_write);
assign ap_return_57 = ~(ap_const_lv288_0_57 ^ lut_out_63_V_write);
assign ap_return_58 = ~(ap_const_lv288_0_58 ^ lut_out_63_V_write);
assign ap_return_59 = ~(ap_const_lv288_0_59 ^ lut_out_63_V_write);
assign ap_return_60 = ~(ap_const_lv288_0_60 ^ lut_out_63_V_write);
assign ap_return_61 = ~(ap_const_lv288_0_61 ^ lut_out_63_V_write);
assign ap_return_62 = ~(ap_const_lv288_0_62 ^ lut_out_63_V_write);
assign ap_return_63 = ~(ap_const_lv288_0_63 ^ lut_out_63_V_write);
endmodule