`timescale 1 ns / 1 ps

module XNORARRAY_b0 (
        lut_out_63_V_write,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63);

parameter    ap_const_lv288_0_0 = 288'h400002000262008000D000010220908A445A001085122041100800200400604000042031;
parameter    ap_const_lv288_0_1 = 288'h8009001C5A000F005A881508A008220402008E2020809588005420048044800000160880;
parameter    ap_const_lv288_0_2 = 288'h2000012000034C02A201508008000010200000100000980000000040002004800000002;
parameter    ap_const_lv288_0_3 = 288'h100A4210D403509E84042808000153A8D018104E26000008A00026084988201050;
parameter    ap_const_lv288_0_4 = 288'h28280080000020810806C4C0000A124082000042880001458519100002080280040080;
parameter    ap_const_lv288_0_5 = 288'h800100024017010201210058002000100280200003002400902002026080868000002042;
parameter    ap_const_lv288_0_6 = 288'h8941802610604E800050800130800D421E1080C040034800240135080402B60000040302;
parameter    ap_const_lv288_0_7 = 288'hC4C80081002B685414A0D890C05500111461801C80E08044440041030110017031488A0;
parameter    ap_const_lv288_0_8 = 288'hC540201050110959281421414008120A0000100001149103294000C92803240800C00208;
parameter    ap_const_lv288_0_9 = 288'h20910690048B191286C30081429C008245039001454280811000408104030092098;
parameter    ap_const_lv288_0_10 = 288'h45B805294011001222020000029C008000030074002518100C5048048514004431001008;
parameter    ap_const_lv288_0_11 = 288'hA8400016A89808001BB8C080001000508030982042000D21380800001000800208032E06;
parameter    ap_const_lv288_0_12 = 288'h40401054C002002080000708412400004000806218400480040300151021400114A14281;
parameter    ap_const_lv288_0_13 = 288'h80404421020200050204C0041002402400020000000E000802508004411000C0040004D4;
parameter    ap_const_lv288_0_14 = 288'h280480C220440C25490CC4858021D4608150D000915458A4000B2034401A000590200406;
parameter    ap_const_lv288_0_15 = 288'h44100001000004C00200049504414431060020D306480420040380100090002101020001;
parameter    ap_const_lv288_0_16 = 288'h2380014042808008005E60280100810000402880400260CC0000C0A00004114022014659;
parameter    ap_const_lv288_0_17 = 288'h464012000000004270892889802A1184300400C0008040804A728720072AA80208D100;
parameter    ap_const_lv288_0_18 = 288'h10058020150005400000900043001A400000260000100008009000840000000820200110;
parameter    ap_const_lv288_0_19 = 288'hE5540801018000858000324000100081008080409441104000704C306441100091084002;
parameter    ap_const_lv288_0_20 = 288'h2440C810246000802008100400E00840000082C01040420004A100C0010202118808820;
parameter    ap_const_lv288_0_21 = 288'h1A0A9E820210D000110A4204180264008240438813420000180C20400010E0011B504884;
parameter    ap_const_lv288_0_22 = 288'h341A84E8C1088020F680084104100420008089201330021922104F988110D5344240849;
parameter    ap_const_lv288_0_23 = 288'h25880E80F000002000A5C518114900580C08017C01A80000215983380A0816600003B88A;
parameter    ap_const_lv288_0_24 = 288'h15B83988053383A050309400D0207B006200013006800D9420009120004900004810432C;
parameter    ap_const_lv288_0_25 = 288'h2A4D2A7000200002284426102A09065208100200234D322338084720184A6080A00A7006;
parameter    ap_const_lv288_0_26 = 288'h4206CCA94302008610020016858000050300004A080488044940084802000C0400027600;
parameter    ap_const_lv288_0_27 = 288'h1001012320106420272810002A600B1C34808100200810B048220010401002000028000;
parameter    ap_const_lv288_0_28 = 288'hA10C0440004004002400804024253400000800300010320003000004092180040280;
parameter    ap_const_lv288_0_29 = 288'h45E05344C082D00691688BC41D4840188A00068112301031284A303050014002320141C0;
parameter    ap_const_lv288_0_30 = 288'h2D8828840F80D80A90023500000620302860820128101A4800200100040204101144600;
parameter    ap_const_lv288_0_31 = 288'h280000221060800146840800100240091002008002446800800840091008002800020454;
parameter    ap_const_lv288_0_32 = 288'h4900802800008C0002D80320000C3A42C00420040200900021832242010512F522908083;
parameter    ap_const_lv288_0_33 = 288'h220006420222002F004200122A0100580A000084044A840104001300400100004000040A;
parameter    ap_const_lv288_0_34 = 288'h10004C41000002088800608000004CC00021001001018810104C400100208011C2888932;
parameter    ap_const_lv288_0_35 = 288'hD0004C2000160684804C4400474681084B10096108440815A04010002400080004081284;
parameter    ap_const_lv288_0_36 = 288'h40080420320000130092881120000001023388210202000000000099012280090002800B;
parameter    ap_const_lv288_0_37 = 288'h9901E086000016C6A8F8868A22202408340100C2000807008581112044049822088510A0;
parameter    ap_const_lv288_0_38 = 288'h400B04040840E24120214142000020000000000A280A0900020030A042801400A002042;
parameter    ap_const_lv288_0_39 = 288'h5D443A020003004A41090160080C028050101404801528E20048110A4A09140650087048;
parameter    ap_const_lv288_0_40 = 288'hC04208000000800C4440508040640000004800302C00518000850502A40085B00C005;
parameter    ap_const_lv288_0_41 = 288'h8010820686000100C43800004000900012880080104040462000480200D621104C7421;
parameter    ap_const_lv288_0_42 = 288'h49484216880901101E2000581545358424028340118007CA8CDA0098B502030508006100;
parameter    ap_const_lv288_0_43 = 288'h88C04A052A4000110001000311062241081000420040200100029680000A240208030231;
parameter    ap_const_lv288_0_44 = 288'h200004602020205800600099040802500440120000098218220806D1010836038200013;
parameter    ap_const_lv288_0_45 = 288'h80012002200102080000400802B10131000000A03821A25D1441230D5C4C0300C40C0008;
parameter    ap_const_lv288_0_46 = 288'hC0820040C08030083105000408416000490021082C904020100310410009000040931;
parameter    ap_const_lv288_0_47 = 288'h4142000000810002034010100AC00003005000240200010210000A048302008645C4EA0;
parameter    ap_const_lv288_0_48 = 288'h2284C802222008C300800801400E0814A00008A120130141081000840400082084129000;
parameter    ap_const_lv288_0_49 = 288'h13880002A8081208400410080210001820A020509008748080B200080045401094006000;
parameter    ap_const_lv288_0_50 = 288'hA000004004200108A001323012C9AE012004000100002801048000B11903002B04C10004;
parameter    ap_const_lv288_0_51 = 288'h10000A000609000700402061600048400009504624002200800B4402840D48440E0;
parameter    ap_const_lv288_0_52 = 288'h508A0320C022112404201A02000344001000400080850844080040041100518C040423C5;
parameter    ap_const_lv288_0_53 = 288'hB02910820901028E89010802112800222000000202000001C1D408801A00808000068820;
parameter    ap_const_lv288_0_54 = 288'h200401950420820400002014288000250E2481B00010151045020042000006040200030;
parameter    ap_const_lv288_0_55 = 288'h82404004022042000A0106018A40000009F0801008800089B10F424458A1CC0150860424;
parameter    ap_const_lv288_0_56 = 288'h4A0840004040008300142020810C04020100000100028040BC00100514010041000C001;
parameter    ap_const_lv288_0_57 = 288'h404060810100184A2002420048620011010209065004232001724C0100000029C00816;
parameter    ap_const_lv288_0_58 = 288'h20204A300420001020100000A0208102AA0020B02202008118768138280D02203C1008F;
parameter    ap_const_lv288_0_59 = 288'h880A014500008001051001900208A00101444400C20011209A0A81010205804104206825;
parameter    ap_const_lv288_0_60 = 288'h148020602080200001A280A81881A064008182010222400A40800A011000011028008000;
parameter    ap_const_lv288_0_61 = 288'h20600918000041300010002804000318C40A0232051000400471000E410A046AA812C00;
parameter    ap_const_lv288_0_62 = 288'h730480100088509410204000340C480024D000C001608108417B408C81817050014DF02;
parameter    ap_const_lv288_0_63 = 288'h800400278014A0341100268140200A48000001C0800046806492243640192001E8401284;
parameter    ap_const_lv288_1_0 = 288'h180408580110100AD9091402800200201100002112809A80490708007020100050001002;
parameter    ap_const_lv288_1_1 = 288'h83480210000000080500004083004008047000A80052016280000000A12482400014040;
parameter    ap_const_lv288_1_2 = 288'h3D1E220148084801900200058954104288010102840442300504081205048B1005000440;
parameter    ap_const_lv288_1_3 = 288'h4BE390270000240124230008B311A11002041228008001004040511AB108A52400006A00;
parameter    ap_const_lv288_1_4 = 288'h220184201580030304548101118081010B4089400052284000000000000092B006080462;
parameter    ap_const_lv288_1_5 = 288'h61C40C820082005008888005342C085880100500818498C4CC290200142485280288900;
parameter    ap_const_lv288_1_6 = 288'h46BE0011001B913401253058020400A4210838080420A40901E248300020400831326080;
parameter    ap_const_lv288_1_7 = 288'h200010024000001A08012000200001580080000000012400200001000028892000000008;
parameter    ap_const_lv288_1_8 = 288'h28E4222824A6600C1CA1C840912C4100416E900180344809002C834101880101117E101;
parameter    ap_const_lv288_1_9 = 288'h210000440000008100080400C48408100240888106408B004210402D0872800902160825;
parameter    ap_const_lv288_1_10 = 288'hB00002420000000100804183A0200E400050460001008040100032521021021000B40600;
parameter    ap_const_lv288_1_11 = 288'h2060921110105A080010008272058094004440100096050C21148AD4025611047200051;
parameter    ap_const_lv288_1_12 = 288'h2805080100C9C800004400200A008482104000000413280931109A2063082E022A120C04;
parameter    ap_const_lv288_1_13 = 288'h441130C0301122C00010180024688AC21088AC4602008001212506122004130000021001;
parameter    ap_const_lv288_1_14 = 288'h52005008400030020030000180801012420001224890208AD4484008000020000010300;
parameter    ap_const_lv288_1_15 = 288'h11E5806C0812802801100002890820400880C0040000900A1A0810001808620200040850;
parameter    ap_const_lv288_1_16 = 288'h458249100202C944B80811184006A1C01128400200C8900204B22050020241041008180;
parameter    ap_const_lv288_1_17 = 288'hA929BC805930142D880060511257C06810CE080212D60013100405185020410404B00800;
parameter    ap_const_lv288_1_18 = 288'h82082080084000800B04282600010010110481400A02AE24204692102A6D249101944865;
parameter    ap_const_lv288_1_19 = 288'h1002860800101F60043880093803A40200005000010A810000008004080800C000308820;
parameter    ap_const_lv288_1_20 = 288'h100200208091143102062732B8196020780E1100A80328C8B00868232044A94845A0292;
parameter    ap_const_lv288_1_21 = 288'h258000005D8028420000012800C110405480206200000400020000082080004004033108;
parameter    ap_const_lv288_1_22 = 288'h4840411008600504006800148045A0DA22200407004F212494A430020009200000800A6;
parameter    ap_const_lv288_1_23 = 288'h20340838828BBB00108222002820C1B28E800011B4BB988224068010C00C85040475;
parameter    ap_const_lv288_1_24 = 288'h8A4042060800680402072001098600339000804010041041100222420032C02400000012;
parameter    ap_const_lv288_1_25 = 288'h4532800C0412802854A2104C14020000200EC8E410300D148001A8012005082300210610;
parameter    ap_const_lv288_1_26 = 288'hC113106108000208AB881A00811080000400024B16066401002E321802222A1087C0982;
parameter    ap_const_lv288_1_27 = 288'h18040A6400B24804990420AD710060480020E28001000204410082100800001280184210;
parameter    ap_const_lv288_1_28 = 288'h99880003089AC19B620D8860462CD0988148109150045E0380141070E8F1640009208441;
parameter    ap_const_lv288_1_29 = 288'h102401000800010000200202070023A0002089020800000042023021800080000A;
parameter    ap_const_lv288_1_30 = 288'h240252206800C025800202952190C08102084001402032538A18014041800D0403007;
parameter    ap_const_lv288_1_31 = 288'h44212500240000180040444001259E0020040B060C000322444501220C44100624F09020;
parameter    ap_const_lv288_1_32 = 288'h400400480950022C00158C4049204B108001021010046300620440008180402850C6440;
parameter    ap_const_lv288_1_33 = 288'h406689AC40900800008D73C40016C600000D0100280142000005402400444021012428A0;
parameter    ap_const_lv288_1_34 = 288'h63942092A4A1310006D48050001030002400302420402041000120000851000808001400;
parameter    ap_const_lv288_1_35 = 288'hE14000A1501895A051001C2089154402009401E9302D48843A024611054017220002450;
parameter    ap_const_lv288_1_36 = 288'h410A20A84ED080820040488100033026480200A01105748C10091020400004040583390;
parameter    ap_const_lv288_1_37 = 288'h20C04010080092001017011C002406300020820443000206002A214A018205120022400;
parameter    ap_const_lv288_1_38 = 288'h8908048005120001400800010318D4A008420440080802085C4484306112D41191120101;
parameter    ap_const_lv288_1_39 = 288'h820040800A0484A00A0240002000400106028888006000118084480000B20021070000A1;
parameter    ap_const_lv288_1_40 = 288'h362208A360038F00B30014020A220AC00A5425EA09019F0842120032004061220042632;
parameter    ap_const_lv288_1_41 = 288'h63A010C1148245C81018200120014420009521802000401090683110015000402A08910;
parameter    ap_const_lv288_1_42 = 288'hB21800025200004052800100024030400558000A1200204104862202404802D0040C51;
parameter    ap_const_lv288_1_43 = 288'h64180500448807004BF200E428000014200412008DA88540040100000420001867C81002;
parameter    ap_const_lv288_1_44 = 288'h24D220804905018208A01822440411980110004C024000822C4F00100005600004400800;
parameter    ap_const_lv288_1_45 = 288'h54BE448909A620B5842C8380090430064240C80A00000020801000C00000004200000400;
parameter    ap_const_lv288_1_46 = 288'h53400450000310884808060502000BA88110002821000002311800086100020420409280;
parameter    ap_const_lv288_1_47 = 288'h930A0450520003159801063042000645042000313201A60302024009108204111A028004;
parameter    ap_const_lv288_1_48 = 288'h44200248C11A800CC9023140035022014200940009084408020400432000001510040204;
parameter    ap_const_lv288_1_49 = 288'h2004AC284012000104F20080514014200204060100428910004C71823000000002028C20;
parameter    ap_const_lv288_1_50 = 288'h48400C3508505C020F7E410F010001001030804C1A0942804200A800A000225073025382;
parameter    ap_const_lv288_1_51 = 288'h23454C00200112944800012810C140911840060100120109081023010300070B02028003;
parameter    ap_const_lv288_1_52 = 288'hA845009320048003290100010A6090004B010611081000002260165200010A7208008008;
parameter    ap_const_lv288_1_53 = 288'h4284892100A0C410001405000012C21803444635404E8400220A204A2490764214306210;
parameter    ap_const_lv288_1_54 = 288'h315002000021040A81246052180040D8080802004640060A5A2008408800F4852902A2C7;
parameter    ap_const_lv288_1_55 = 288'h49F9152E410304C641A90266431B433020F5123D040A54004208109020C11A20B219918;
parameter    ap_const_lv288_1_56 = 288'h1483053000C4204B49800840003800003C119064415909001000320100128022729C0;
parameter    ap_const_lv288_1_57 = 288'h4B59903049488000058210009A58062020400000009000441140011000A200110090000;
parameter    ap_const_lv288_1_58 = 288'hC01B14C80148002445C8FA1945010208100102008CA0BE0200880040810041080040040;
parameter    ap_const_lv288_1_59 = 288'h2B008205081481222CD4023401010C08018034225B244850055084229504D8889481000;
parameter    ap_const_lv288_1_60 = 288'h420800000138081782154E554248140000100084908430C00002004864020006C0042475;
parameter    ap_const_lv288_1_61 = 288'h912110084140030841008B0C1C114204110841000008C8000210008A0208410800000004;
parameter    ap_const_lv288_1_62 = 288'h90802002000002000204B003A0000B020000005020000280100002100080000000802009;
parameter    ap_const_lv288_1_63 = 288'h44021000000010062601908014301200206040141149118130082810940800804948840;


input  [287:0] lut_out_63_V_write;
output  [287:0] ap_return_0;
output  [287:0] ap_return_1;
output  [287:0] ap_return_2;
output  [287:0] ap_return_3;
output  [287:0] ap_return_4;
output  [287:0] ap_return_5;
output  [287:0] ap_return_6;
output  [287:0] ap_return_7;
output  [287:0] ap_return_8;
output  [287:0] ap_return_9;
output  [287:0] ap_return_10;
output  [287:0] ap_return_11;
output  [287:0] ap_return_12;
output  [287:0] ap_return_13;
output  [287:0] ap_return_14;
output  [287:0] ap_return_15;
output  [287:0] ap_return_16;
output  [287:0] ap_return_17;
output  [287:0] ap_return_18;
output  [287:0] ap_return_19;
output  [287:0] ap_return_20;
output  [287:0] ap_return_21;
output  [287:0] ap_return_22;
output  [287:0] ap_return_23;
output  [287:0] ap_return_24;
output  [287:0] ap_return_25;
output  [287:0] ap_return_26;
output  [287:0] ap_return_27;
output  [287:0] ap_return_28;
output  [287:0] ap_return_29;
output  [287:0] ap_return_30;
output  [287:0] ap_return_31;
output  [287:0] ap_return_32;
output  [287:0] ap_return_33;
output  [287:0] ap_return_34;
output  [287:0] ap_return_35;
output  [287:0] ap_return_36;
output  [287:0] ap_return_37;
output  [287:0] ap_return_38;
output  [287:0] ap_return_39;
output  [287:0] ap_return_40;
output  [287:0] ap_return_41;
output  [287:0] ap_return_42;
output  [287:0] ap_return_43;
output  [287:0] ap_return_44;
output  [287:0] ap_return_45;
output  [287:0] ap_return_46;
output  [287:0] ap_return_47;
output  [287:0] ap_return_48;
output  [287:0] ap_return_49;
output  [287:0] ap_return_50;
output  [287:0] ap_return_51;
output  [287:0] ap_return_52;
output  [287:0] ap_return_53;
output  [287:0] ap_return_54;
output  [287:0] ap_return_55;
output  [287:0] ap_return_56;
output  [287:0] ap_return_57;
output  [287:0] ap_return_58;
output  [287:0] ap_return_59;
output  [287:0] ap_return_60;
output  [287:0] ap_return_61;
output  [287:0] ap_return_62;
output  [287:0] ap_return_63;
assign ap_return_0 = (ap_const_lv288_0_0 & lut_out_63_V_write) | (ap_const_lv288_1_0 & ~lut_out_63_V_write);
assign ap_return_1 = (ap_const_lv288_0_1 & lut_out_63_V_write) | (ap_const_lv288_1_1 & ~lut_out_63_V_write);
assign ap_return_2 = (ap_const_lv288_0_2 & lut_out_63_V_write) | (ap_const_lv288_1_2 & ~lut_out_63_V_write);
assign ap_return_3 = (ap_const_lv288_0_3 & lut_out_63_V_write) | (ap_const_lv288_1_3 & ~lut_out_63_V_write);
assign ap_return_4 = (ap_const_lv288_0_4 & lut_out_63_V_write) | (ap_const_lv288_1_4 & ~lut_out_63_V_write);
assign ap_return_5 = (ap_const_lv288_0_5 & lut_out_63_V_write) | (ap_const_lv288_1_5 & ~lut_out_63_V_write);
assign ap_return_6 = (ap_const_lv288_0_6 & lut_out_63_V_write) | (ap_const_lv288_1_6 & ~lut_out_63_V_write);
assign ap_return_7 = (ap_const_lv288_0_7 & lut_out_63_V_write) | (ap_const_lv288_1_7 & ~lut_out_63_V_write);
assign ap_return_8 = (ap_const_lv288_0_8 & lut_out_63_V_write) | (ap_const_lv288_1_8 & ~lut_out_63_V_write);
assign ap_return_9 = (ap_const_lv288_0_9 & lut_out_63_V_write) | (ap_const_lv288_1_9 & ~lut_out_63_V_write);
assign ap_return_10 = (ap_const_lv288_0_10 & lut_out_63_V_write) | (ap_const_lv288_1_10 & ~lut_out_63_V_write);
assign ap_return_11 = (ap_const_lv288_0_11 & lut_out_63_V_write) | (ap_const_lv288_1_11 & ~lut_out_63_V_write);
assign ap_return_12 = (ap_const_lv288_0_12 & lut_out_63_V_write) | (ap_const_lv288_1_12 & ~lut_out_63_V_write);
assign ap_return_13 = (ap_const_lv288_0_13 & lut_out_63_V_write) | (ap_const_lv288_1_13 & ~lut_out_63_V_write);
assign ap_return_14 = (ap_const_lv288_0_14 & lut_out_63_V_write) | (ap_const_lv288_1_14 & ~lut_out_63_V_write);
assign ap_return_15 = (ap_const_lv288_0_15 & lut_out_63_V_write) | (ap_const_lv288_1_15 & ~lut_out_63_V_write);
assign ap_return_16 = (ap_const_lv288_0_16 & lut_out_63_V_write) | (ap_const_lv288_1_16 & ~lut_out_63_V_write);
assign ap_return_17 = (ap_const_lv288_0_17 & lut_out_63_V_write) | (ap_const_lv288_1_17 & ~lut_out_63_V_write);
assign ap_return_18 = (ap_const_lv288_0_18 & lut_out_63_V_write) | (ap_const_lv288_1_18 & ~lut_out_63_V_write);
assign ap_return_19 = (ap_const_lv288_0_19 & lut_out_63_V_write) | (ap_const_lv288_1_19 & ~lut_out_63_V_write);
assign ap_return_20 = (ap_const_lv288_0_20 & lut_out_63_V_write) | (ap_const_lv288_1_20 & ~lut_out_63_V_write);
assign ap_return_21 = (ap_const_lv288_0_21 & lut_out_63_V_write) | (ap_const_lv288_1_21 & ~lut_out_63_V_write);
assign ap_return_22 = (ap_const_lv288_0_22 & lut_out_63_V_write) | (ap_const_lv288_1_22 & ~lut_out_63_V_write);
assign ap_return_23 = (ap_const_lv288_0_23 & lut_out_63_V_write) | (ap_const_lv288_1_23 & ~lut_out_63_V_write);
assign ap_return_24 = (ap_const_lv288_0_24 & lut_out_63_V_write) | (ap_const_lv288_1_24 & ~lut_out_63_V_write);
assign ap_return_25 = (ap_const_lv288_0_25 & lut_out_63_V_write) | (ap_const_lv288_1_25 & ~lut_out_63_V_write);
assign ap_return_26 = (ap_const_lv288_0_26 & lut_out_63_V_write) | (ap_const_lv288_1_26 & ~lut_out_63_V_write);
assign ap_return_27 = (ap_const_lv288_0_27 & lut_out_63_V_write) | (ap_const_lv288_1_27 & ~lut_out_63_V_write);
assign ap_return_28 = (ap_const_lv288_0_28 & lut_out_63_V_write) | (ap_const_lv288_1_28 & ~lut_out_63_V_write);
assign ap_return_29 = (ap_const_lv288_0_29 & lut_out_63_V_write) | (ap_const_lv288_1_29 & ~lut_out_63_V_write);
assign ap_return_30 = (ap_const_lv288_0_30 & lut_out_63_V_write) | (ap_const_lv288_1_30 & ~lut_out_63_V_write);
assign ap_return_31 = (ap_const_lv288_0_31 & lut_out_63_V_write) | (ap_const_lv288_1_31 & ~lut_out_63_V_write);
assign ap_return_32 = (ap_const_lv288_0_32 & lut_out_63_V_write) | (ap_const_lv288_1_32 & ~lut_out_63_V_write);
assign ap_return_33 = (ap_const_lv288_0_33 & lut_out_63_V_write) | (ap_const_lv288_1_33 & ~lut_out_63_V_write);
assign ap_return_34 = (ap_const_lv288_0_34 & lut_out_63_V_write) | (ap_const_lv288_1_34 & ~lut_out_63_V_write);
assign ap_return_35 = (ap_const_lv288_0_35 & lut_out_63_V_write) | (ap_const_lv288_1_35 & ~lut_out_63_V_write);
assign ap_return_36 = (ap_const_lv288_0_36 & lut_out_63_V_write) | (ap_const_lv288_1_36 & ~lut_out_63_V_write);
assign ap_return_37 = (ap_const_lv288_0_37 & lut_out_63_V_write) | (ap_const_lv288_1_37 & ~lut_out_63_V_write);
assign ap_return_38 = (ap_const_lv288_0_38 & lut_out_63_V_write) | (ap_const_lv288_1_38 & ~lut_out_63_V_write);
assign ap_return_39 = (ap_const_lv288_0_39 & lut_out_63_V_write) | (ap_const_lv288_1_39 & ~lut_out_63_V_write);
assign ap_return_40 = (ap_const_lv288_0_40 & lut_out_63_V_write) | (ap_const_lv288_1_40 & ~lut_out_63_V_write);
assign ap_return_41 = (ap_const_lv288_0_41 & lut_out_63_V_write) | (ap_const_lv288_1_41 & ~lut_out_63_V_write);
assign ap_return_42 = (ap_const_lv288_0_42 & lut_out_63_V_write) | (ap_const_lv288_1_42 & ~lut_out_63_V_write);
assign ap_return_43 = (ap_const_lv288_0_43 & lut_out_63_V_write) | (ap_const_lv288_1_43 & ~lut_out_63_V_write);
assign ap_return_44 = (ap_const_lv288_0_44 & lut_out_63_V_write) | (ap_const_lv288_1_44 & ~lut_out_63_V_write);
assign ap_return_45 = (ap_const_lv288_0_45 & lut_out_63_V_write) | (ap_const_lv288_1_45 & ~lut_out_63_V_write);
assign ap_return_46 = (ap_const_lv288_0_46 & lut_out_63_V_write) | (ap_const_lv288_1_46 & ~lut_out_63_V_write);
assign ap_return_47 = (ap_const_lv288_0_47 & lut_out_63_V_write) | (ap_const_lv288_1_47 & ~lut_out_63_V_write);
assign ap_return_48 = (ap_const_lv288_0_48 & lut_out_63_V_write) | (ap_const_lv288_1_48 & ~lut_out_63_V_write);
assign ap_return_49 = (ap_const_lv288_0_49 & lut_out_63_V_write) | (ap_const_lv288_1_49 & ~lut_out_63_V_write);
assign ap_return_50 = (ap_const_lv288_0_50 & lut_out_63_V_write) | (ap_const_lv288_1_50 & ~lut_out_63_V_write);
assign ap_return_51 = (ap_const_lv288_0_51 & lut_out_63_V_write) | (ap_const_lv288_1_51 & ~lut_out_63_V_write);
assign ap_return_52 = (ap_const_lv288_0_52 & lut_out_63_V_write) | (ap_const_lv288_1_52 & ~lut_out_63_V_write);
assign ap_return_53 = (ap_const_lv288_0_53 & lut_out_63_V_write) | (ap_const_lv288_1_53 & ~lut_out_63_V_write);
assign ap_return_54 = (ap_const_lv288_0_54 & lut_out_63_V_write) | (ap_const_lv288_1_54 & ~lut_out_63_V_write);
assign ap_return_55 = (ap_const_lv288_0_55 & lut_out_63_V_write) | (ap_const_lv288_1_55 & ~lut_out_63_V_write);
assign ap_return_56 = (ap_const_lv288_0_56 & lut_out_63_V_write) | (ap_const_lv288_1_56 & ~lut_out_63_V_write);
assign ap_return_57 = (ap_const_lv288_0_57 & lut_out_63_V_write) | (ap_const_lv288_1_57 & ~lut_out_63_V_write);
assign ap_return_58 = (ap_const_lv288_0_58 & lut_out_63_V_write) | (ap_const_lv288_1_58 & ~lut_out_63_V_write);
assign ap_return_59 = (ap_const_lv288_0_59 & lut_out_63_V_write) | (ap_const_lv288_1_59 & ~lut_out_63_V_write);
assign ap_return_60 = (ap_const_lv288_0_60 & lut_out_63_V_write) | (ap_const_lv288_1_60 & ~lut_out_63_V_write);
assign ap_return_61 = (ap_const_lv288_0_61 & lut_out_63_V_write) | (ap_const_lv288_1_61 & ~lut_out_63_V_write);
assign ap_return_62 = (ap_const_lv288_0_62 & lut_out_63_V_write) | (ap_const_lv288_1_62 & ~lut_out_63_V_write);
assign ap_return_63 = (ap_const_lv288_0_63 & lut_out_63_V_write) | (ap_const_lv288_1_63 & ~lut_out_63_V_write);
endmodule